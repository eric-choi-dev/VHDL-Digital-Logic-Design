library verilog;
use verilog.vl_types.all;
entity Jcounter_vlg_vec_tst is
end Jcounter_vlg_vec_tst;
